// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8

module c499 (keyinput2,N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input [15:0] keyinput2;
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;

output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723;

wire N724_OBFUS,N725_OBFUS,N726_OBFUS,N727_OBFUS,N728_OBFUS,N729_OBFUS,N730_OBFUS,N731_OBFUS,N732_OBFUS,N733_OBFUS,
       N734_OBFUS,N735_OBFUS,N736_OBFUS,N737_OBFUS,N738_OBFUS,N739_OBFUS,N740_OBFUS,N741_OBFUS,N742_OBFUS,N743_OBFUS,
       N744_OBFUS,N745_OBFUS,N746_OBFUS,N747_OBFUS,N748_OBFUS,N749_OBFUS,N750_OBFUS,N751_OBFUS,N752_OBFUS,N753_OBFUS,
       N754_OBFUS,N755_OBFUS;

xor XOR2_1 (N250, N1, N5);
xor XOR2_2 (N251, N9, N13);
xor XOR2_3 (N252, N17, N21);
xor XOR2_4 (N253, N25, N29);
xor XOR2_5 (N254, N33, N37);
xor XOR2_6 (N255, N41, N45);
xor XOR2_7 (N256, N49, N53);
xor XOR2_8 (N257, N57, N61);
xor XOR2_9 (N258, N65, N69);
xor XOR2_10 (N259, N73, N77);
xor XOR2_11 (N260, N81, N85);
xor XOR2_12 (N261, N89, N93);
xor XOR2_13 (N262, N97, N101);
xor XOR2_14 (N263, N105, N109);
xor XOR2_15 (N264, N113, N117);
xor XOR2_16 (N265, N121, N125);
and AND2_17 (N266, N129, N137);
and AND2_18 (N267, N130, N137);
and AND2_19 (N268, N131, N137);
and AND2_20 (N269, N132, N137);
and AND2_21 (N270, N133, N137);
and AND2_22 (N271, N134, N137);
and AND2_23 (N272, N135, N137);
and AND2_24 (N273, N136, N137);
xor XOR2_25 (N274, N1, N17);
xor XOR2_26 (N275, N33, N49);
xor XOR2_27 (N276, N5, N21);
xor XOR2_28 (N277, N37, N53);
xor XOR2_29 (N278, N9, N25);
xor XOR2_30 (N279, N41, N57);
xor XOR2_31 (N280, N13, N29);
xor XOR2_32 (N281, N45, N61);
xor XOR2_33 (N282, N65, N81);
xor XOR2_34 (N283, N97, N113);
xor XOR2_35 (N284, N69, N85);
xor XOR2_36 (N285, N101, N117);
xor XOR2_37 (N286, N73, N89);
xor XOR2_38 (N287, N105, N121);
xor XOR2_39 (N288, N77, N93);
xor XOR2_40 (N289, N109, N125);
xor XOR2_41 (N290, N250, N251);
xor XOR2_42 (N293, N252, N253);
xor XOR2_43 (N296, N254, N255);
xor XOR2_44 (N299, N256, N257);
xor XOR2_45 (N302, N258, N259);
xor XOR2_46 (N305, N260, N261);
xor XOR2_47 (N308, N262, N263);
xor XOR2_48 (N311, N264, N265);
xor XOR2_49 (N314, N274, N275);
xor XOR2_50 (N315, N276, N277);
xor XOR2_51 (N316, N278, N279);
xor XOR2_52 (N317, N280, N281);
xor XOR2_53 (N318, N282, N283);
xor XOR2_54 (N319, N284, N285);
xor XOR2_55 (N320, N286, N287);
xor XOR2_56 (N321, N288, N289);
xor XOR2_57 (N338, N290, N293);
xor XOR2_58 (N339, N296, N299);
xor XOR2_59 (N340, N290, N296);
xor XOR2_60 (N341, N293, N299);
xor XOR2_61 (N342, N302, N305);
xor XOR2_62 (N343, N308, N311);
xor XOR2_63 (N344, N302, N308);
xor XOR2_64 (N345, N305, N311);
xor XOR2_65 (N346, N266, N342);
xor XOR2_66 (N347, N267, N343);
xor XOR2_67 (N348, N268, N344);
xor XOR2_68 (N349, N269, N345);
xor XOR2_69 (N350, N270, N338);
xor XOR2_70 (N351, N271, N339);
xor XOR2_71 (N352, N272, N340);
xor XOR2_72 (N353, N273, N341);
xor XOR2_73 (N354, N314, N346);
xor XOR2_74 (N367, N315, N347);
xor XOR2_75 (N380, N316, N348);
xor XOR2_76 (N393, N317, N349);
xor XOR2_77 (N406, N318, N350);
xor XOR2_78 (N419, N319, N351);
xor XOR2_79 (N432, N320, N352);
xor XOR2_80 (N445, N321, N353);
not NOT1_81 (N554, N354);
not NOT1_82 (N555, N367);
not NOT1_83 (N556, N380);
not NOT1_84 (N557, N354);
not NOT1_85 (N558, N367);
not NOT1_86 (N559, N393);
not NOT1_87 (N560, N354);
not NOT1_88 (N561, N380);
not NOT1_89 (N562, N393);
not NOT1_90 (N563, N367);
not NOT1_91 (N564, N380);
not NOT1_92 (N565, N393);
not NOT1_93 (N566, N419);
not NOT1_94 (N567, N445);
not NOT1_95 (N568, N419);
not NOT1_96 (N569, N432);
not NOT1_97 (N570, N406);
not NOT1_98 (N571, N445);
not NOT1_99 (N572, N406);
not NOT1_100 (N573, N432);
not NOT1_101 (N574, N406);
not NOT1_102 (N575, N419);
not NOT1_103 (N576, N432);
not NOT1_104 (N577, N406);
not NOT1_105 (N578, N419);
not NOT1_106 (N579, N445);
not NOT1_107 (N580, N406);
not NOT1_108 (N581, N432);
not NOT1_109 (N582, N445);
not NOT1_110 (N583, N419);
not NOT1_111 (N584, N432);
not NOT1_112 (N585, N445);
not NOT1_113 (N586, N367);
not NOT1_114 (N587, N393);
not NOT1_115 (N588, N367);
not NOT1_116 (N589, N380);
not NOT1_117 (N590, N354);
not NOT1_118 (N591, N393);
not NOT1_119 (N592, N354);
not NOT1_120 (N593, N380);
and AND4_121 (N594, N554, N555, N556, N393);
and AND4_122 (N595, N557, N558, N380, N559);
and AND4_123 (N596, N560, N367, N561, N562);
and AND4_124 (N597, N354, N563, N564, N565);
and AND4_125 (N598, N574, N575, N576, N445);
and AND4_126 (N599, N577, N578, N432, N579);
and AND4_127 (N600, N580, N419, N581, N582);
and AND4_128 (N601, N406, N583, N584, N585);
or OR4_129 (N602, N594, N595, N596, N597);
or OR4_130 (N607, N598, N599, N600, N601);
and AND5_131 (N620, N406, N566, N432, N567, N602);
and AND5_132 (N625, N406, N568, N569, N445, N602);
and AND5_133 (N630, N570, N419, N432, N571, N602);
and AND5_134 (N635, N572, N419, N573, N445, N602);
and AND5_135 (N640, N354, N586, N380, N587, N607);
and AND5_136 (N645, N354, N588, N589, N393, N607);
and AND5_137 (N650, N590, N367, N380, N591, N607);
and AND5_138 (N655, N592, N367, N593, N393, N607);
and AND2_139 (N692, N354, N620);
and AND2_140 (N693, N367, N620);
and AND2_141 (N694, N380, N620);
and AND2_142 (N695, N393, N620);
and AND2_143 (N696, N354, N625);
and AND2_144 (N697, N367, N625);
and AND2_145 (N698, N380, N625);
and AND2_146 (N699, N393, N625);
and AND2_147 (N700, N354, N630);
and AND2_148 (N701, N367, N630);
and AND2_149 (N702, N380, N630);
and AND2_150 (N703, N393, N630);
and AND2_151 (N704, N354, N635);
and AND2_152 (N705, N367, N635);
and AND2_153 (N706, N380, N635);
and AND2_154 (N707, N393, N635);
and AND2_155 (N708, N406, N640);
and AND2_156 (N709, N419, N640);
and AND2_157 (N710, N432, N640);
and AND2_158 (N711, N445, N640);
and AND2_159 (N712, N406, N645);
and AND2_160 (N713, N419, N645);
and AND2_161 (N714, N432, N645);
and AND2_162 (N715, N445, N645);
and AND2_163 (N716, N406, N650);
and AND2_164 (N717, N419, N650);
and AND2_165 (N718, N432, N650);
and AND2_166 (N719, N445, N650);
and AND2_167 (N720, N406, N655);
and AND2_168 (N721, N419, N655);
and AND2_169 (N722, N432, N655);
and AND2_170 (N723, N445, N655);
xor XOR2_171 (N724_OBFUS, N1, N692);
xor XOR2_171_OBFUS (N724, N724_OBFUS, keyinput2[0]);

xor XOR2_172 (N725_OBFUS, N5, N693);
xnor XOR2_172_OBFUS (N725, N725_OBFUS, keyinput2[1]);

xor XOR2_173 (N726_OBFUS, N9, N694);
xnor XOR2_173_OBFUS (N726, N726_OBFUS, keyinput2[2]);

xor XOR2_174 (N727_OBFUS, N13, N695);
xnor XOR2_174_OBFUS (N727, N727_OBFUS, keyinput2[4]);

xor XOR2_175 (N728_OBFUS, N17, N696);
xor XOR2_175_OBFUS (N728, N728_OBFUS, keyinput2[7]);

xor XOR2_176 (N729_OBFUS, N21, N697);
xnor XOR2_176_OBFUS (N729, N729_OBFUS, keyinput2[3]);

xor XOR2_177 (N730_OBFUS, N25, N698);
xor XOR2_177_OBFUS (N730, N730_OBFUS, keyinput2[5]);

xor XOR2_178 (N731_OBFUS, N29, N699);
xnor XOR2_178_OBFUS (N731, N731_OBFUS, keyinput2[6]);

xor XOR2_179 (N732_OBFUS, N33, N700);
xor XOR2_179_OBFUS (N732, N732_OBFUS, keyinput2[9]);

xor XOR2_180 (N733_OBFUS, N37, N701);
xnor XOR2_180_OBFUS (N733, N733_OBFUS, keyinput2[8]);

xor XOR2_181 (N734_OBFUS, N41, N702);
xor XOR2_181_OBFUS (N734, N734_OBFUS, keyinput2[10]);

xor XOR2_182 (N735_OBFUS, N45, N703);
xnor XOR2_182_OBFUS (N735, N735_OBFUS, keyinput2[11]); 

xor XOR2_183 (N736_OBFUS, N49, N704);
xnor XOR2_183_OBFUS (N736, N736_OBFUS, keyinput2[12]);

xor XOR2_184 (N737_OBFUS, N53, N705);
xnor XOR2_184_OBFUS (N737, N737_OBFUS, keyinput2[13]);

xor XOR2_185 (N738_OBFUS, N57, N706);
xnor XOR2_185_OBFUS (N738, N738_OBFUS, keyinput2[14]);

xor XOR2_186 (N739_OBFUS, N61, N707);
xor XOR2_186_OBFUS (N739, N739_OBFUS, keyinput2[15]);

xor XOR2_187 (N740, N65, N708);
xor XOR2_188 (N741, N69, N709);
xor XOR2_189 (N742, N73, N710);
xor XOR2_190 (N743, N77, N711);
xor XOR2_191 (N744, N81, N712);
xor XOR2_192 (N745, N85, N713);
xor XOR2_193 (N746, N89, N714);
xor XOR2_194 (N747, N93, N715);
xor XOR2_195 (N748, N97, N716);
xor XOR2_196 (N749, N101, N717);
xor XOR2_197 (N750, N105, N718);
xor XOR2_198 (N751, N109, N719);
xor XOR2_199 (N752, N113, N720);
xor XOR2_200 (N753, N117, N721);
xor XOR2_201 (N754, N121, N722);
xor XOR2_202 (N755, N125, N723);

endmodule
